module C_XOR(
input A,
input B,
output OUT
);

  assign OUT = A^B;
endmodule
